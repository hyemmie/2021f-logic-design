`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:15:52 10/14/2021 
// Design Name: 
// Module Name:    dLatchAndFlipFlop 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dLatchAndFlipFlop(
    input D,
    input CLK,
    output Qlatch,
    output Qflipflop
    );
	 
	 wire temp1;
	 wire temp2;
	 
	 dLatch dl(D, CLK, Qlatch, temp1);
	 dFlipFlop dff(D, CLK, Qflipflop, temp2);


endmodule
